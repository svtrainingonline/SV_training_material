module shree_ganesha();

initial
  begin
    $display ("Shree Ganesha");
  end
endmodule
